/*
* Copyright (c) 2025. All rights reserved.
* Created by dulat, 10/17/25
*/

module top #(
    parameter [7:0] WIDTH = 8'h0
) (
    input  wire [7:0] in,
    output wire [7:0] out
);

    assign out = in;

endmodule
